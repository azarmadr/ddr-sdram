initial begin : test

cke     <=  1'b0;
cs_n    <=  1'b1;
ras_n   <=  1'b1;
cas_n   <=  1'b1;
we_n    <=  1'b1;
ba      <=  {BA_BITS{1'bz}};
a       <=  {ADDR_BITS{1'bz}};
dq_en   <=  1'b0;
dqs_en  <=  1'b0;
cke     <=  1'b1;
power_up;
$display("Powerup complete");
precharge('h00000000, 1);
nop(trp);
load_mode('h1, 'h00002000);
nop(tmrd-1);
load_mode('h0, 'h0000013A);
nop(tmrd-1);
precharge('h00000000, 1);
nop(trp);
refresh;
nop(trfc);
refresh;
nop(trfc);
load_mode('h0, 'h0000003A);
nop(tmrd-1);
nop('h000000C8);
activate('h00000000, 'h00000000);
nop(trcd-1);
write('h00000000, 'h00000000, 1, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30003000, 32'h20002000, 32'h10001000, 32'h0});
nop(BL/2+twr);
activate('h00000001, 'h00000000);
nop(trcd-1);
write('h00000001, 'h00000000, 1, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30013001, 32'h20012001, 32'h10011001, 32'h10001});
nop(BL/2+twr);
activate('h00000002, 'h00000000);
nop(trcd-1);
write('h00000002, 'h00000000, 1, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30023002, 32'h20022002, 32'h10021002, 32'h20002});
nop(BL/2+twr);
activate('h00000003, 'h00000000);
nop(trcd-1);
write('h00000003, 'h00000000, 1, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30033003, 32'h20032003, 32'h10031003, 32'h30003});
nop(BL/2+twr);
activate('h00000000, 'h00000000);
nop(trrd-1);
activate('h00000001, 'h00000000);
nop(trrd-1);
activate('h00000002, 'h00000000);
nop(trrd-1);
activate('h00000003, 'h00000000);
read('h00000000, 'h00000000, 1);
nop(BL/2-1);
read('h00000001, 'h00000000, 1);
nop(BL/2-1);
read('h00000002, 'h00000000, 1);
nop(BL/2-1);
read('h00000003, 'h00000000, 1);
nop(BL/2+twr-2);
activate('h00000001, 'h00000000);
nop(trrd-1);
activate('h00000000, 'h00000000);
nop(trcd-1);
$display("%m At time %t: WRITE Burst", $time);write('h00000000, 'h00000004, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30403040, 32'h20402040, 32'h10401040, 32'h400040});
nop(BL/2+4);
$display("%m At time %t: Consecutive WRITE to WRITE", $time);write('h00000000, 'h00000008, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h30803080, 32'h20802080, 32'h10801080, 32'h800080});
nop(BL/2-1);
write('h00000000, 'h0000000C, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h31203120, 32'h21202120, 32'h11201120, 32'h1200120});
nop(BL/2-1);
$display("%m At time %t: Nonconsecutive WRITE to WRITE", $time);write('h00000000, 'h00000010, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h31603160, 32'h21602160, 32'h11601160, 32'h1600160});
nop(BL/2+4);
write('h00000000, 'h00000014, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h32003200, 32'h22002200, 32'h12001200, 32'h2000200});
nop(BL/2+twr+4);
$display("%m At time %t: Random WRITE Cycles", $time);write('h00000000, 'h00000018, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h32403240, 32'h22402240, 32'h12401240, 32'h2400240});
nop(BL/2-1);
write('h00000000, 'h0000001C, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h32803280, 32'h22802280, 32'h12801280, 32'h2800280});
nop(BL/2-1);
write('h00000000, 'h00000020, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h33203320, 32'h23202320, 32'h13201320, 32'h3200320});
nop(BL/2-1);
write('h00000000, 'h00000024, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h33603360, 32'h23602360, 32'h13601360, 32'h3600360});
nop(BL/2-1);
$display("%m At time %t: WRITE to READ - Uninterrupting", $time);write('h00000000, 'h00000028, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h34003400, 32'h24002400, 32'h14001400, 32'h4000400});
nop(BL/2+1);
read('h00000000, 'h00000028, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Interrupting", $time);write('h00000000, 'h0000002C, 0, { 4'h1, 4'h1, 4'h0, 4'h0}, { 32'h34403440, 32'h24402440, 32'h14401440, 32'h4400440});
nop(BL/2+1);
read('h00000000, 'h0000002C, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Odd Number of Data, Interrupting", $time);write('h00000000, 'h00000030, 0, { 4'h1, 4'h1, 4'h1, 4'h0}, { 32'h34803480, 32'h24802480, 32'h14801480, 32'h4800480});
nop(BL/2+1);
read('h00000000, 'h00000030, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to PRECHARGE - Uninterrupting", $time);write('h00000000, 'h00000034, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h35203520, 32'h25202520, 32'h15201520, 32'h5200520});
nop(BL/2+twr);
precharge('h00000000, 0);
nop(trp-1);
$display("%m At time %t: WRITE with AUTO PRECHARGE", $time);activate('h00000000, 'h00000000);
nop(trcd-1);
write('h00000000, 'h00000040, 1, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h36603660, 32'h26602660, 32'h16601660, 32'h6600660});
nop(BL/2+twr+trp);
activate('h00000000, 'h00000000);
nop(trcd-1);
$display("%m At time %t: READ Burst", $time);read('h00000000, 'h00000000, 0);
nop(BL/2-1);
$display("%m At time %t: Consecutive READ Bursts", $time);read('h00000000, 'h00000004, 0);
nop(BL/2-2);
read('h00000000, 'h00000008, 0);
nop(BL/2-1);
$display("%m At time %t: Nonconsecutive READ Bursts", $time);read('h00000000, 'h0000000C, 0);
nop(BL/2);
read('h00000000, 'h00000010, 0);
nop(BL/2);
$display("%m At time %t: Random READ Accesses", $time);read('h00000000, 'h00000014, 0);
read('h00000000, 'h00000018, 0);
read('h00000000, 'h0000001C, 0);
read('h00000000, 'h00000020, 0);
nop(BL/2);
$display("%m At time %t: Terminating a READ Burst", $time);read('h00000000, 'h00000024, 0);
burst_term;
nop(BL/2-2);
$display("%m At time %t: READ to WRITE", $time);read('h00000000, 'h00000028, 0);
burst_term;
nop(CL);
write('h00000000, 'h0000002C, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'h34C034C0, 32'h24C024C0, 32'h14C014C0, 32'h4C004C0});
nop(BL/2+1);
$display("%m At time %t: READ to PRECHARGE", $time);read('h00000000, 'h00000030, 0);
nop('h00000001);
precharge('h00000000, 0);
nop(trp-1);
$display("%m At time %t: READ with AUTO PRECHARGE", $time);activate('h00000000, 'h00000000);
nop(trcd-1);
read('h00000000, 'h00000034, 1);
nop(CL+BL/2+twr);
$display("%m At time %t: WRITE to READ - Mask byte 0 of Burst 0", $time);activate('h00000000, 'h00000000);
nop(trcd-1);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h1}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 1 of Burst 0", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h2}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 2 of Burst 0", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h4}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 3 of Burst 0", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h8}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 0 of Burst 1", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h1, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 1 of Burst 1", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h2, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 2 of Burst 1", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h4, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 3 of Burst 1", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h8, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 0 of Burst 2", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h1, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 1 of Burst 2", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h2, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 2 of Burst 2", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h4, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 3 of Burst 2", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h0, 4'h8, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 0 of Burst 3", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h1, 4'h0, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 1 of Burst 3", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h2, 4'h0, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 2 of Burst 3", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h4, 4'h0, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 0);
nop(CL+BL/2-1);
$display("%m At time %t: WRITE to READ - Mask byte 3 of Burst 3", $time);write('h00000000, 'h00000064, 0, { 4'h0, 4'h0, 4'h0, 4'h0}, { 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
nop(BL/2);
write('h00000000, 'h00000064, 0, { 4'h8, 4'h0, 4'h0, 4'h0}, { 32'h33333333, 32'h22222222, 32'h11111111, 32'h0});
nop(BL/2+1);
read('h00000000, 'h00000064, 1);
nop(CL+BL/2-1);
test_done = 1;
end

